/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module SC_TRANSICION_NIVEL (
	//////////// OUTPUTS //////////
	DATA_FIXED_INITREGPOINT_7_OutBUS,
	DATA_FIXED_INITREGPOINT_6_OutBUS,
	DATA_FIXED_INITREGPOINT_5_OutBUS,
	DATA_FIXED_INITREGPOINT_4_OutBUS,
	DATA_FIXED_INITREGPOINT_3_OutBUS,
	DATA_FIXED_INITREGPOINT_2_OutBUS,
	DATA_FIXED_INITREGPOINT_1_OutBUS,
	DATA_FIXED_INITREGPOINT_0_OutBUS,
	
	DATA_FIXED_INITREGBACKG_7_OutBUS,
	DATA_FIXED_INITREGBACKG_6_OutBUS,
	DATA_FIXED_INITREGBACKG_5_OutBUS,
	DATA_FIXED_INITREGBACKG_4_OutBUS,
	DATA_FIXED_INITREGBACKG_3_OutBUS,
	DATA_FIXED_INITREGBACKG_2_OutBUS,
	DATA_FIXED_INITREGBACKG_1_OutBUS,
	DATA_FIXED_INITREGBACKG_0_OutBUS,
	//////////// INPUTS //////////
	SC_RegNIVEL_CLOCK_50,
	SC_RegNIVEL_RESET_InHigh,
	SC_RegNIVEL_clear_InLow, 
	SC_RegNIVEL_load_InLow, 
	
	DATA_FIXED_INITREGPOINT_7_InBUS,
	DATA_FIXED_INITREGPOINT_6_InBUS,
	DATA_FIXED_INITREGPOINT_5_InBUS,
	DATA_FIXED_INITREGPOINT_4_InBUS
	DATA_FIXED_INITREGPOINT_3_InBUS,
	DATA_FIXED_INITREGPOINT_2_InBUS,
	DATA_FIXED_INITREGPOINT_1_InBUS,
	DATA_FIXED_INITREGPOINT_0_InBUS,
	
	DATA_FIXED_INITREGBACKG_7_InBUS,
	DATA_FIXED_INITREGBACKG_6_InBUS,
	DATA_FIXED_INITREGBACKG_5_InBUS,
	DATA_FIXED_INITREGBACKG_4_InBUS,
	DATA_FIXED_INITREGBACKG_3_InBUS,
	DATA_FIXED_INITREGBACKG_2_InBUS,
	DATA_FIXED_INITREGBACKG_1_InBUS,
	DATA_FIXED_INITREGBACKG_0_InBUS,
	
	STATEMACHINE_MAIN_transition_InBUS


);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output[8-1:0] DATA_FIXED_INITREGPOINT_7_InBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_7_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_6_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_5_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_4_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_3_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_2_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_1_OutBUS;
output[8-1:0] DATA_FIXED_INITREGPOINT_0_OutBUS;
	
output[8-1:0] DATA_FIXED_INITREGBACKG_7_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_6_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_5_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_4_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_3_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_2_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_1_OutBUS;
output[8-1:0] DATA_FIXED_INITREGBACKG_0_OutBUS;


input		SC_RegNIVEL_CLOCK_50;
input		SC_RegNIVEL_RESET_InHigh;
input		SC_RegNIVEL_clear_InLow;
input		SC_RegNIVEL_load_InLow;	


input[8-1:0] DATA_FIXED_INITREGPOINT_7_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_6_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_5_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_4_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_3_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_2_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_1_InBUS;
input[8-1:0] DATA_FIXED_INITREGPOINT_0_InBUS;

input[8-1:0] DATA_FIXED_INITREGBACKG_7_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_6_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_5_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_4_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_3_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_2_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_1_InBUS,
input[8-1:0] DATA_FIXED_INITREGBACKG_0_InBUS


//=======================================================
//  REG/WIRE declarations
//=======================================================
reg [8-1:0] RegNIVEL_Register;
reg [8-1:0] RegNIVEL_Signal;
//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
always @(*) 
begin

	if (STATEMACHINE_MAIN_transition_cwire == 3b'001) begin

		 DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_0 = 8'b00000000;

		 DATA_FIXED_INITREGBACKG_7 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_6 = 8'b00011000;
		 DATA_FIXED_INITREGBACKG_5 = 8'b00111000;
		 DATA_FIXED_INITREGBACKG_4 = 8'b00011000;
		 DATA_FIXED_INITREGBACKG_3 = 8'b00011000;
		 DATA_FIXED_INITREGBACKG_2 = 8'b00011000;
		 DATA_FIXED_INITREGBACKG_1 = 8'b00111100;
		 DATA_FIXED_INITREGBACKG_0 = 8'b00000000;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3b'010) begin

		 DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_FIXED_INITREGBACKG_7 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_6 = 8'b00111000;
		 DATA_FIXED_INITREGBACKG_5 = 8'b01000100;
		 DATA_FIXED_INITREGBACKG_4 = 8'b00001000;
		 DATA_FIXED_INITREGBACKG_3 = 8'b00010000;
		 DATA_FIXED_INITREGBACKG_2 = 8'b00100000;
		 DATA_FIXED_INITREGBACKG_1 = 8'b01111100;
		 DATA_FIXED_INITREGBACKG_0 = 8'b00000000;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3b'011) begin

		 DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_FIXED_INITREGBACKG_7 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_6 = 8'b01111100;
		 DATA_FIXED_INITREGBACKG_5 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_4 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_3 = 8'b01111100;
		 DATA_FIXED_INITREGBACKG_2 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_1 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_0 = 8'b01111110;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3b'100) begin

		 DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_FIXED_INITREGBACKG_7 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_6 = 8'b01000010;
		 DATA_FIXED_INITREGBACKG_5 = 8'b01000010;
		 DATA_FIXED_INITREGBACKG_4 = 8'b01000010;
		 DATA_FIXED_INITREGBACKG_3 = 8'b01111010;
		 DATA_FIXED_INITREGBACKG_2 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_1 = 8'b00000010;
		 DATA_FIXED_INITREGBACKG_0 = 8'b00000000;
		 end
		
	else begin

		 DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
		 DATA_FIXED_INITREGPOINT_0 = 8'b00010000;
		 
		
		 DATA_FIXED_INITREGBACKG_7 = 8'b11100000;
		 DATA_FIXED_INITREGBACKG_6 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_5 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_4 = 8'b11100000;
		 DATA_FIXED_INITREGBACKG_3 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_2 = 8'b11100000;
		 DATA_FIXED_INITREGBACKG_1 = 8'b00000000;
		 DATA_FIXED_INITREGBACKG_0 = 8'b00000000;
		 end
	 
	 end 
//STATE REGISTER: SEQUENTIAL
always @(posedge SC_RegNIVEL_CLOCK_50, posedge SC_RegNIVEL_RESET_InHigh)
begin
	if (SC_RegNIVEL_RESET_InHigh == 1'b1)
		RegNIVEL_Register <= 0;
	else
		RegNIVEL_Register <= RegNIVEL_Signal;
end
//=======================================================
//  Outputs
//=======================================================
//OUTPUT LOGIC: COMBINATIONAL
assign SC_RegNIVEL_data_OutBUS = RegNIVEL_Register;

endmodule