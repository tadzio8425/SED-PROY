



module CC_SET_FIXED_TRANSITIONS (
	
		/////// OUTPUTS ////////////////////////
		 DATA_TRANSITION_INITREGPOINT_7,
		 DATA_TRANSITION_INITREGPOINT_6,
		 DATA_TRANSITION_INITREGPOINT_5,
		 DATA_TRANSITION_INITREGPOINT_4,
		 DATA_TRANSITION_INITREGPOINT_3,
		 DATA_TRANSITION_INITREGPOINT_2,
		 DATA_TRANSITION_INITREGPOINT_1,
		 DATA_TRANSITION_INITREGPOINT_0,

		 DATA_TRANSITION_INITREGBACKG_7,
		 DATA_TRANSITION_INITREGBACKG_6,
		 DATA_TRANSITION_INITREGBACKG_5,
		 DATA_TRANSITION_INITREGBACKG_4,
		 DATA_TRANSITION_INITREGBACKG_3,
		 DATA_TRANSITION_INITREGBACKG_2,
		 DATA_TRANSITION_INITREGBACKG_1,
		 DATA_TRANSITION_INITREGBACKG_0,
		 
		///////// INPUTS ///////////////////////

		 STATEMACHINE_MAIN_transition_cwire
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output reg  [8-1:0]   DATA_TRANSITION_INITREGPOINT_7;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_6;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_5;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_4;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_3;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_2;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_1;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGPOINT_0;

output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_7;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_6;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_5;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_4;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_3;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_2;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_1;
output reg	[8-1:0]	 DATA_TRANSITION_INITREGBACKG_0;

input STATEMACHINE_MAIN_transition_cwire;

//=======================================================
//  REG/WIRE declarations
//=======================================================



//=======================================================
//  Structural coding
//=======================================================
always @(*) 
begin

	if (STATEMACHINE_MAIN_transition_cwire == 3'b001) begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00000000;

		 DATA_TRANSITION_INITREGBACKG_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b00111000;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b00111100;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b00000000;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3'b010) begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_TRANSITION_INITREGBACKG_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b00111000;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b01000100;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b00001000;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b00010000;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b00100000;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b01111100;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b00000000;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3'b011) begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_TRANSITION_INITREGBACKG_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b01111100;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b01111100;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b01111110;
		 end
		 
		 
	else if (STATEMACHINE_MAIN_transition_cwire == 3'b100) begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_TRANSITION_INITREGBACKG_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b01000010;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b01000010;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b01000010;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b01111010;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b00000010;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b00000000;
		
		 end
		 
	
	else if (STATEMACHINE_MAIN_transition_cwire == 3'b101) begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00000000;
		 
		 
		 //////////// POS INICIAL FONDO / OBSTACULOS /////
		 DATA_TRANSITION_INITREGBACKG_7 = 8'b11111111;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b01111110;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b01111110;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b01111110;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b00011000;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b00111100;
		
		 end
		 		 
		
	else begin

		 DATA_TRANSITION_INITREGPOINT_7 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_4 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_2 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGPOINT_0 = 8'b00010000;
		 
		
		 DATA_TRANSITION_INITREGBACKG_7 = 8'b11011011;
		 DATA_TRANSITION_INITREGBACKG_6 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_5 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_4 = 8'b11100000;
		 DATA_TRANSITION_INITREGBACKG_3 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_2 = 8'b11100000;
		 DATA_TRANSITION_INITREGBACKG_1 = 8'b00000000;
		 DATA_TRANSITION_INITREGBACKG_0 = 8'b00000000;
		 end
	 
	 end 
endmodule
