//=======================================================
//  MODULE Definition
//=======================================================
module CC_COLLISION_DETECTOR #(parameter COLLISION_DETECTOR_DATAWIDTH=8)(
	

	CC_COLLISION_DETECTOR_OutLow,
		/////////// INPUTS //////////
	CC_COLLISION_DETECTOR_BACK_InBUS_u0,
	CC_COLLISION_DETECTOR_BACK_InBUS_u1,
	CC_COLLISION_DETECTOR_BACK_InBUS_u2,
	CC_COLLISION_DETECTOR_BACK_InBUS_u3,
	CC_COLLISION_DETECTOR_BACK_InBUS_u4,
	CC_COLLISION_DETECTOR_BACK_InBUS_u5,
	CC_COLLISION_DETECTOR_BACK_InBUS_u6,
	CC_COLLISION_DETECTOR_BACK_InBUS_u7,
	
	CC_COLLISION_DETECTOR_POINT_InBUS_u0,
	CC_COLLISION_DETECTOR_POINT_InBUS_u1,
	CC_COLLISION_DETECTOR_POINT_InBUS_u2,
	CC_COLLISION_DETECTOR_POINT_InBUS_u3,
	CC_COLLISION_DETECTOR_POINT_InBUS_u4,
	CC_COLLISION_DETECTOR_POINT_InBUS_u5,
	CC_COLLISION_DETECTOR_POINT_InBUS_u6,
	CC_COLLISION_DETECTOR_POINT_InBUS_u7
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output	reg CC_COLLISION_DETECTOR_OutLow;


input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u0;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u1;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u2;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u3;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u4;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u5;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u6;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_BACK_InBUS_u7;
	
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u0;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u1;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u2;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u3;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u4;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u5;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u6;
input 	[COLLISION_DETECTOR_DATAWIDTH-1:0]	CC_COLLISION_DETECTOR_POINT_InBUS_u7;


//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
always @(*)
begin
	if( (CC_COLLISION_DETECTOR_POINT_InBUS_u7 & CC_COLLISION_DETECTOR_BACK_InBUS_u7) != 8'b00000000 ||
	    (CC_COLLISION_DETECTOR_POINT_InBUS_u6 & CC_COLLISION_DETECTOR_BACK_InBUS_u6) != 8'b00000000 ||
	    (CC_COLLISION_DETECTOR_POINT_InBUS_u5 & CC_COLLISION_DETECTOR_BACK_InBUS_u5) != 8'b00000000 ||
		 (CC_COLLISION_DETECTOR_POINT_InBUS_u4 & CC_COLLISION_DETECTOR_BACK_InBUS_u4) != 8'b00000000 ||
		 (CC_COLLISION_DETECTOR_POINT_InBUS_u3 & CC_COLLISION_DETECTOR_BACK_InBUS_u3) != 8'b00000000 ||
		 (CC_COLLISION_DETECTOR_POINT_InBUS_u2 & CC_COLLISION_DETECTOR_BACK_InBUS_u2) != 8'b00000000 ||
		 (CC_COLLISION_DETECTOR_POINT_InBUS_u1 & CC_COLLISION_DETECTOR_BACK_InBUS_u1) != 8'b00000000 ||
		 (CC_COLLISION_DETECTOR_POINT_InBUS_u0 & CC_COLLISION_DETECTOR_BACK_InBUS_u0) != 8'b00000000 )
	
		CC_COLLISION_DETECTOR_OutLow = 1'b0;
	else 
		CC_COLLISION_DETECTOR_OutLow = 1'b1;
end

endmodule


